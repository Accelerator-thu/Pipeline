module Control (OpCode,
                Funct);
    input [5:0] OpCode, Funct;
    
endmodule
