module Pipeline (
    clk,
    reset,
    out
);
    input clk;
    input reset;
    output out;

    
endmodule