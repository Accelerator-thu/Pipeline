module Forward(clk,
               reset,
               );
    
endmodule
