module RegEXMEM ();
    
endmodule
